`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Engineer: Ryan Bride (For Northeastern UN LAB) 
// Create Date: 08/02/2023 01:55:36 PM
// Module Name: MAC
// Project Name: 40Gb/s (And 100Gb/s Ethernet Core) 
// Description: Top File For the MAC  
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//      First Version Exist to Talk to RS layer For timing Reasons with
//      PCS, RS layer is not The standard they defined in the EEE manual
//      But achieves the same thing 
//////////////////////////////////////////////////////////////////////////////////
module MAC(

    );
    
    
    
endmodule
